package top_package;

    
    parameter CHIP_ADDR     = 8'hCD;
    parameter SCCB_CLKDIV   = 12'd125;


endpackage