package top_package;

    // ov7670 sccb parameters //
    parameter CHIP_ADDR     = 8'hCD;
    parameter SCCB_CLKDIV   = 12'd125;
    // ov7670 sccb parameters //


endpackage