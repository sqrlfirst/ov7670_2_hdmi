module im_compression_tb;

    localparam in_width = ;

    logic [639:0][479:0][2:0][7:0]        pic_batman;



    initial begin
        pic_batman = $readmem(batman.mem)
    end




endmodule 
